// Joash Shankar, Ming He, Nikhil Pillai
// ECE 5760 Final Project Spring 2024
// Blackjack
// DE1_SoC_Computer.v

module DE1_SoC_Computer (
	////////////////////////////////////
	// FPGA Pins
	////////////////////////////////////

	// Clock pins
	CLOCK_50,
	CLOCK2_50,
	CLOCK3_50,
	CLOCK4_50,

	// ADC
	ADC_CS_N,
	ADC_DIN,
	ADC_DOUT,
	ADC_SCLK,

	// Audio
	AUD_ADCDAT,
	AUD_ADCLRCK,
	AUD_BCLK,
	AUD_DACDAT,
	AUD_DACLRCK,
	AUD_XCK,

	// SDRAM
	DRAM_ADDR,
	DRAM_BA,
	DRAM_CAS_N,
	DRAM_CKE,
	DRAM_CLK,
	DRAM_CS_N,
	DRAM_DQ,
	DRAM_LDQM,
	DRAM_RAS_N,
	DRAM_UDQM,
	DRAM_WE_N,

	// I2C Bus for Configuration of the Audio and Video-In Chips
	FPGA_I2C_SCLK,
	FPGA_I2C_SDAT,

	// 40-Pin Headers
	GPIO_0,
	GPIO_1,
	
	// Seven Segment Displays
	HEX0,
	HEX1,
	HEX2,
	HEX3,
	HEX4,
	HEX5,

	// IR
	IRDA_RXD,
	IRDA_TXD,

	// Pushbuttons
	KEY,

	// LEDs
	LEDR,

	// PS2 Ports
	PS2_CLK,
	PS2_DAT,
	
	PS2_CLK2,
	PS2_DAT2,

	// Slider Switches
	SW,

	// Video-In
	TD_CLK27,
	TD_DATA,
	TD_HS,
	TD_RESET_N,
	TD_VS,

	// VGA
	VGA_B,
	VGA_BLANK_N,
	VGA_CLK,
	VGA_G,
	VGA_HS,
	VGA_R,
	VGA_SYNC_N,
	VGA_VS,

	////////////////////////////////////
	// HPS Pins
	////////////////////////////////////
	
	// DDR3 SDRAM
	HPS_DDR3_ADDR,
	HPS_DDR3_BA,
	HPS_DDR3_CAS_N,
	HPS_DDR3_CKE,
	HPS_DDR3_CK_N,
	HPS_DDR3_CK_P,
	HPS_DDR3_CS_N,
	HPS_DDR3_DM,
	HPS_DDR3_DQ,
	HPS_DDR3_DQS_N,
	HPS_DDR3_DQS_P,
	HPS_DDR3_ODT,
	HPS_DDR3_RAS_N,
	HPS_DDR3_RESET_N,
	HPS_DDR3_RZQ,
	HPS_DDR3_WE_N,

	// Ethernet
	HPS_ENET_GTX_CLK,
	HPS_ENET_INT_N,
	HPS_ENET_MDC,
	HPS_ENET_MDIO,
	HPS_ENET_RX_CLK,
	HPS_ENET_RX_DATA,
	HPS_ENET_RX_DV,
	HPS_ENET_TX_DATA,
	HPS_ENET_TX_EN,

	// Flash
	HPS_FLASH_DATA,
	HPS_FLASH_DCLK,
	HPS_FLASH_NCSO,

	// Accelerometer
	HPS_GSENSOR_INT,
		
	// General Purpose I/O
	HPS_GPIO,
		
	// I2C
	HPS_I2C_CONTROL,
	HPS_I2C1_SCLK,
	HPS_I2C1_SDAT,
	HPS_I2C2_SCLK,
	HPS_I2C2_SDAT,

	// Pushbutton
	HPS_KEY,

	// LED
	HPS_LED,
		
	// SD Card
	HPS_SD_CLK,
	HPS_SD_CMD,
	HPS_SD_DATA,

	// SPI
	HPS_SPIM_CLK,
	HPS_SPIM_MISO,
	HPS_SPIM_MOSI,
	HPS_SPIM_SS,

	// UART
	HPS_UART_RX,
	HPS_UART_TX,

	// USB
	HPS_CONV_USB_N,
	HPS_USB_CLKOUT,
	HPS_USB_DATA,
	HPS_USB_DIR,
	HPS_USB_NXT,
	HPS_USB_STP,
);

//=======================================================
//  PARAMETER declarations
//=======================================================


//=======================================================
//  PORT declarations
//=======================================================

////////////////////////////////////
// FPGA Pins
////////////////////////////////////

// Clock pins
input						CLOCK_50;
input						CLOCK2_50;
input						CLOCK3_50;
input						CLOCK4_50;

// ADC
inout						ADC_CS_N;
output					ADC_DIN;
input						ADC_DOUT;
output					ADC_SCLK;

// Audio
input						AUD_ADCDAT;
inout						AUD_ADCLRCK;
inout						AUD_BCLK;
output					AUD_DACDAT;
inout						AUD_DACLRCK;
output					AUD_XCK;

// SDRAM
output 		[12: 0]	DRAM_ADDR;
output		[ 1: 0]	DRAM_BA;
output					DRAM_CAS_N;
output					DRAM_CKE;
output					DRAM_CLK;
output					DRAM_CS_N;
inout			[15: 0]	DRAM_DQ;
output					DRAM_LDQM;
output					DRAM_RAS_N;
output					DRAM_UDQM;
output					DRAM_WE_N;

// I2C Bus for Configuration of the Audio and Video-In Chips
output					FPGA_I2C_SCLK;
inout						FPGA_I2C_SDAT;

// 40-pin headers
inout			[35: 0]	GPIO_0;
inout			[35: 0]	GPIO_1;

// Seven Segment Displays
output		[ 6: 0]	HEX0;
output		[ 6: 0]	HEX1;
output		[ 6: 0]	HEX2;
output		[ 6: 0]	HEX3;
output		[ 6: 0]	HEX4;
output		[ 6: 0]	HEX5;

// IR
input						IRDA_RXD;
output					IRDA_TXD;

// Pushbuttons
input			[ 3: 0]	KEY;

// LEDs
output		[ 9: 0]	LEDR;

// PS2 Ports
inout						PS2_CLK;
inout						PS2_DAT;

inout						PS2_CLK2;
inout						PS2_DAT2;

// Slider Switches
input			[ 9: 0]	SW;

// Video-In
input						TD_CLK27;
input			[ 7: 0]	TD_DATA;
input						TD_HS;
output					TD_RESET_N;
input						TD_VS;

// VGA
output		[ 7: 0]	VGA_B;
output					VGA_BLANK_N;
output					VGA_CLK;
output		[ 7: 0]	VGA_G;
output					VGA_HS;
output		[ 7: 0]	VGA_R;
output					VGA_SYNC_N;
output					VGA_VS;



////////////////////////////////////
// HPS Pins
////////////////////////////////////
	
// DDR3 SDRAM
output		[14: 0]	HPS_DDR3_ADDR;
output		[ 2: 0]  HPS_DDR3_BA;
output					HPS_DDR3_CAS_N;
output					HPS_DDR3_CKE;
output					HPS_DDR3_CK_N;
output					HPS_DDR3_CK_P;
output					HPS_DDR3_CS_N;
output		[ 3: 0]	HPS_DDR3_DM;
inout			[31: 0]	HPS_DDR3_DQ;
inout			[ 3: 0]	HPS_DDR3_DQS_N;
inout			[ 3: 0]	HPS_DDR3_DQS_P;
output					HPS_DDR3_ODT;
output					HPS_DDR3_RAS_N;
output					HPS_DDR3_RESET_N;
input						HPS_DDR3_RZQ;
output					HPS_DDR3_WE_N;

// Ethernet
output					HPS_ENET_GTX_CLK;
inout						HPS_ENET_INT_N;
output					HPS_ENET_MDC;
inout						HPS_ENET_MDIO;
input						HPS_ENET_RX_CLK;
input			[ 3: 0]	HPS_ENET_RX_DATA;
input						HPS_ENET_RX_DV;
output		[ 3: 0]	HPS_ENET_TX_DATA;
output					HPS_ENET_TX_EN;

// Flash
inout			[ 3: 0]	HPS_FLASH_DATA;
output					HPS_FLASH_DCLK;
output					HPS_FLASH_NCSO;

// Accelerometer
inout						HPS_GSENSOR_INT;

// General Purpose I/O
inout			[ 1: 0]	HPS_GPIO;

// I2C
inout						HPS_I2C_CONTROL;
inout						HPS_I2C1_SCLK;
inout						HPS_I2C1_SDAT;
inout						HPS_I2C2_SCLK;
inout						HPS_I2C2_SDAT;

// Pushbutton
inout						HPS_KEY;

// LED
inout						HPS_LED;

// SD Card
output					HPS_SD_CLK;
inout						HPS_SD_CMD;
inout			[ 3: 0]	HPS_SD_DATA;

// SPI
output					HPS_SPIM_CLK;
input						HPS_SPIM_MISO;
output					HPS_SPIM_MOSI;
inout						HPS_SPIM_SS;

// UART
input						HPS_UART_RX;
output					HPS_UART_TX;

// USB
inout						HPS_CONV_USB_N;
input						HPS_USB_CLKOUT;
inout			[ 7: 0]	HPS_USB_DATA;
input						HPS_USB_DIR;
input						HPS_USB_NXT;
output					HPS_USB_STP;

//=======================================================
//  REG/WIRE declarations
//=======================================================

wire			[31: 0]	hex3_hex0;
//wire			[15: 0]	hex5_hex4;

assign HEX0 = hex3_hex0[ 3: 0]; // hex3_hex0[ 6: 0]; 
assign HEX1 = hex3_hex0[7: 4];
assign HEX2 = hex3_hex0[11:8];
assign HEX3 = hex3_hex0[15:12];
assign HEX4 = hex3_hex0[19:16];
assign HEX5 = hex3_hex0[23:20];

//HexDigit Digit0(HEX0, hex3_hex0[3:0]);
//HexDigit Digit1(HEX1, hex3_hex0[7:4]);
//HexDigit Digit2(HEX2, hex3_hex0[11:8]);
//HexDigit Digit3(HEX3, hex3_hex0[15:12]);

// VGA clock and reset lines
wire vga_pll_lock ;
wire vga_pll ;
reg  vga_reset ;
assign hex3_hex = max_time;
// M10k memory control and data
wire 		[7:0] 	M10k_out [15:0];
wire 		[7:0] 	write_data [15:0];
wire 		[18:0] 	write_address [15:0];
reg 		[18:0] 	read_address ;
wire 					write_enable [15:0];
wire	         write_enable_2;
//Second M10k block
wire 		[7:0] 	M10k_out_2 ;
wire 		[7:0] 	write_data_2;// stores color data
wire 		[18:0] 	write_address_2 ;
wire 		[18:0] 	read_address_2 ;

// M10k memory clock
wire 					M10k_pll /*synthesis keep */;
wire 					M10k_pll_locked ;

// Memory writing control registers
reg 		[7:0] 	arbiter_state ;
wire 		[9:0] 	x_coord ;
wire 		[9:0] 	y_coord ;
wire 		[9:0] 	x_coord_2 ;
wire 		[9:0] 	y_coord_2;

// initial values for x and y 
reg [9:0] init_x [1:0];
reg [9:0] init_y [1:0];

// Wires for connecting VGA driver to memory
wire 		[9:0]		next_x ;
wire 		[9:0] 	next_y ;

// wires for ci, cr, and max_iter
reg signed [26:0] ci, cr, ci_2, cr_2;
wire [11:0] counter [15:0];
wire [11:0] counter_2;
wire [11:0] max_iterations;
assign max_iterations = 12'd1000;

wire calc_done [15:0];
wire calc_done_2;

wire [26:0] unit_step_size_cr, step_size_cr, step_size_ci;

assign unit_step_size_cr = {4'b0000, 23'b00000001001100110011001} >> pio_zoom_cr_external_connection_export[5:0]; 
assign step_size_cr = ({4'b0000, 23'b00000010011001100110010}) >> pio_zoom_cr_external_connection_export[5:0];
assign step_size_ci = {4'b0000, 23'b00000001000100010001000} >> pio_zoom_ci_external_connection_export[5:0];

//KEY debouncing -> seems not necessary
//key_debouncing state_3(.clk(M10k_pll), .button_in(KEY[3]), .button_state(button_state_3));
//key_debouncing state_2(.clk(M10k_pll), .button_in(KEY[2]), .button_state(button_state_2));
//key_debouncing state_1(.clk(M10k_pll), .button_in(KEY[1]), .button_state(button_state_1));
//wire [1:0] button_state_0;
//key_debouncing state_0(.clk(M10k_pll), .button_in(KEY[0]), .button_state(button_state_0));

// wire for time counter
wire [31:0] counter_external_connection_export;
wire flag_counter;

reg [3:0] itr_counter; // counter loops 16 iterators and keeps the max time to send to HPS
reg [31:0] time_inter_data, max_time; // timer to keep the intermediate time data
reg [15:0] record_flag; 

wire time_flag [15:0];
wire time_flag_2;

wire [31:0] time_counter [15:0];
wire [31:0] time_counter_2;
reg [31:0] t_counter, t_counter_2;

assign counter_external_connection_export = max_time; 

always@(posedge M10k_pll) begin	
	// four buttons to move the graph
	if(pio_reset_external_connection_export[0] || ~KEY[0]) begin
		itr_counter <= 0;
		max_time <= 0;
	end
	else begin
//	if(time_flag[0] && time_flag[1] && time_flag[2] && time_flag[3] && time_flag[4] && time_flag[5] && time_flag[6] && time_flag[7] &&
//		time_flag[8] && time_flag[9] && time_flag[10] && time_flag[11] && time_flag[12] && time_flag[13] && time_flag[14] && time_flag[15] ) begin
		if(time_flag[0]) begin
			record_flag <= record_flag | 16'd1;
		end
		if(time_flag[1]) begin
			record_flag <= record_flag | (16'd1 << 1);
		end
		if(time_flag[2]) begin
			record_flag <= record_flag | (16'd1 << 2);
		end
		if(time_flag[3]) begin
			record_flag <= record_flag | (16'd1 << 3);
		end
		if(time_flag[4]) begin
			record_flag <= record_flag | (16'd1 << 4);
		end
		if(time_flag[5]) begin
			record_flag <= record_flag | (16'd1 << 5);
		end
		if(time_flag[6]) begin
			record_flag <= record_flag | (16'd1 << 6);
		end
		if(time_flag[7]) begin
			record_flag <= record_flag | (16'd1 << 7);
		end
		if(time_flag[8]) begin
			record_flag <= record_flag | (16'd1 << 8);
		end
		if(time_flag[9]) begin
			record_flag <= record_flag | (16'd1 << 9);
		end
		if(time_flag[10]) begin
			record_flag <= record_flag | (16'd1 << 10);
		end
		if(time_flag[11]) begin
			record_flag <= record_flag | (16'd1 << 11);
		end
		if(time_flag[12]) begin
			record_flag <= record_flag | (16'd1 << 12);
		end
		if(time_flag[13]) begin
			record_flag <= record_flag | (16'd1 << 13);
		end
		if(time_flag[14]) begin
			record_flag <= record_flag | (16'd1 << 14);
		end
		if(time_flag[15]) begin
			record_flag <= record_flag | (16'd1 << 15);
		end
				
		itr_counter <= itr_counter + 1;
		case(itr_counter)
        4'd0: time_inter_data = time_counter[0];
        4'd1: time_inter_data = time_counter[1];
        4'd2: time_inter_data = time_counter[2];
        4'd3: time_inter_data = time_counter[3];
        4'd4: time_inter_data = time_counter[4];
        4'd5: time_inter_data = time_counter[5];
        4'd6: time_inter_data = time_counter[6];
        4'd7: time_inter_data = time_counter[7];
        4'd8: time_inter_data = time_counter[8];
        4'd9: time_inter_data = time_counter[9];
        4'd10: time_inter_data = time_counter[10];
        4'd11: time_inter_data = time_counter[11];
        4'd12: time_inter_data = time_counter[12];
        4'd13: time_inter_data = time_counter[13];
        4'd14: time_inter_data = time_counter[14];
        4'd15: time_inter_data = time_counter[15];
		  default time_inter_data = 32'd0 ;
      endcase
	max_time <= (max_time <= time_inter_data) ? time_inter_data : max_time;
	if (itr_counter > 15) begin
		itr_counter <= 0;
	end
	if(&record_flag) begin
		max_time <= 0;
		record_flag <= 0;
	end
	end
end

//assign step_size_x = ({4'b0000, 23'b00000001001100110011001} << 1) >> SW[5:0];
//assign step_every_other_x = ({4'b0000, 23'b00000010011001100110010}) >> SW[5:0];
//assign step_size_x = {4'b0000, 23'b00000001001100110011001}; //3/640
//assign step_size_y = {4'b0000, 23'b00000001000100010001000} >> SW[5:0];
//assign LEDR[0] = (~KEY[3]) ? 1'd1 : 1'd0;
//assign LEDR[1] = (~KEY[0]) ? 1'd1 : 1'd0;

// wires for ci/cr increment/zoom and pio reset
wire [31:0] pio_ci_init_external_connection_export;
wire [31:0] pio_cr_init_external_connection_export;
wire [31:0] pio_zoom_ci_external_connection_export;
wire [31:0] pio_zoom_cr_external_connection_export;
wire [7:0] pio_reset_external_connection_export;

// wire for max iterations
wire [15:0] pio_max_iter_external_connection_export;
 
wire [18:0] calc_address;
assign calc_address = ((19'd_40*next_y) + (next_x >> 4));

wire [7:0] color_in_VGA_inter [15:0];
//assign color_in_VGA = next_x[0] ? M10k_out_2 : M10k_out;

wire [7:0] color_in_VGA;

/*
reg [18:0] mem_block_index ; 
always@(*)
begin
    case(next_x[3:0])
        6'd0: mem_block_index=M10K_out[0];
        6'd1: mem_block_index=1;
        6'd2: mem_block_index=32'd2925946;
        6'd3: mem_block_index=32'd3284755;
        6'd4: mem_block_index=32'd3686513;
        6'd5: mem_block_index=32'd3905735;
        6'd6: mem_block_index=32'd4384445;
        6'd7: mem_block_index=32'd4921316;
        6'd8: mem_block_index=32'd5524401;
        6'd9: mem_block_index=32'd5852787;
        6'd10: mem_block_index=32'd6569510;
        6'd11: mem_block_index=32'd7373921;
        6'd12: mem_block_index=32'd7812366;
        6'd13: mem_block_index=32'd8768891;
        6'd14: mem_block_index=32'd9842633;
        6'd15: mem_block_index=32'd11047908;
        default mem_block_index =32'd0 ;
    endcase
end
*/

genvar i;
generate
	for (i=0; i<16; i=i+1) begin: instBlocks
		mandelbrot MBROT (.clock(M10k_pll),
								.reset(pio_reset_external_connection_export[0] || ~KEY[0]),				
								.x_coord_init(10'd_0+i),
								.y_coord_init(10'd_0),
//								.step_size_cr(step_size_cr),
                        .step_size_cr(unit_step_size_cr << 4),
								.step_size_ci(step_size_ci),
								.c_i_init(pio_ci_init_external_connection_export[26:0]),
								.c_r_init(pio_cr_init_external_connection_export[26:0] + (i * unit_step_size_cr)),
								.max_iter(pio_max_iter_external_connection_export),
								.out(counter[i]),
								.write_en (write_enable[i]),
								.write_addr(write_address[i]),
								.done(calc_done[i]),
								.time_flag(time_flag[i]),
								.time_counter(time_counter[i]));		
		
		M10K_1000_8 pixel_data( .q(M10k_out[i]), // contains pixel color (8 bit) for display
										.d(write_data[i]),
										.write_address(write_address[i]),
										.read_address(calc_address),
										.we(write_enable[i]),
										.clk(M10k_pll));
		
		// assign color_in_VGA_inter[i] = next_x[0] ? M10k_out[0] : M10k_out[1];
		
		color_write color_iter(.clk(M10k_pll), 
										.counter(counter[i]), 
										.max_iterations(pio_max_iter_external_connection_export), 
										.write_data_out(write_data[i]));						
										
	end
endgenerate

//assign color_in_VGA = next_x[0] ? M10k_out[1] : M10k_out[0];
//assign color_in_VGA = color_in_VGA_inter[0];
assign color_in_VGA = M10k_out[next_x[3:0]];
/*
// Instantiate memory
M10K_1000_8 pixel_data( .q(M10k_out), // contains pixel color (8 bit) for display
								.d(write_data),
								.write_address(write_address),
								.read_address(calc_address),
								.we(write_enable),
								.clk(M10k_pll)
);


M10K_1000_8 pixel_data_2( .q(M10k_out_2), // contains pixel color (8 bit) for display
								.d(write_data_2),
								.write_address(write_address_2),
								.read_address(calc_address),
								.we(write_enable_2),
								.clk(M10k_pll)
);
*/

// Instantiate VGA driver					
vga_driver DUT   (	.clock(vga_pll), 
							.reset(pio_reset_external_connection_export[0] || ~KEY[0]),
							.color_in(color_in_VGA),	// Pixel color (8-bit) from memory
							.next_x(next_x),		// This (and next_y) used to specify memory read address
							.next_y(next_y),		// This (and next_x) used to specify memory read address
							.hsync(VGA_HS),
							.vsync(VGA_VS),
							.red(VGA_R),
							.green(VGA_G),
							.blue(VGA_B),
							.sync(VGA_SYNC_N),
							.clk(VGA_CLK),
							.blank(VGA_BLANK_N)
);


/*
// Instantiation of Mandelbrot
    mandelbrot MBROT (.clock(M10k_pll),
            .reset(pio_reset_external_connection_export[0] || ~KEY[0]),				
			   .x_coord_init(10'd_0),
			   .y_coord_init(10'd_0),
				.step_size_cr(step_size_cr),
				.step_size_ci(step_size_ci),
            .c_i_init(pio_ci_init_external_connection_export[26:0]),
				.c_r_init(pio_cr_init_external_connection_export[26:0]),
				//.c_i_init({4'b0001, 23'd0}),
				//.c_r_init({-4'b0010, 23'd0}),
				.max_iter(max_iterations),
				.out(counter),
				.write_en (write_enable),
				.write_addr(write_address),
				.done(calc_done),
				.time_flag(time_flag),
				.time_counter(time_counter)	);
    
	mandelbrot MBROT_2 (.clock(M10k_pll),
            .reset(pio_reset_external_connection_export[0] || ~KEY[0]),
			   .x_coord_init(10'd_1),
			   .y_coord_init(10'd_0),			
				.step_size_cr(step_size_cr),
				.step_size_ci(step_size_ci),
            .c_i_init(pio_ci_init_external_connection_export[26:0]),
				.c_r_init(pio_cr_init_external_connection_export[26:0] + unit_step_size_cr),
				//.c_i_init({4'b0001, 23'd0}),
			   //.c_r_init({4'sb1110, 23'b00000001001100110011001}),
				//.c_r_init({-4'b0010, 23'd0} + ({4'b0000, 23'b00000001001100110011001} >> SW[5:0])),
				.max_iter(max_iterations),
				.out(counter_2),
				.write_en(write_enable_2),
				.write_addr(write_address_2),
				.done(calc_done_2),
				.time_flag(time_flag_2),
				.time_counter(time_counter_2)	);

// Instantiation of color write data
color_write color_iterOne(.clk(M10k_pll), .counter(counter), .max_iterations(max_iterations), .write_data_out(write_data));
color_write color_iterTwo(.clk(M10k_pll), .counter(counter_2), .max_iterations(max_iterations), .write_data_out(write_data_2));
*/
	
//=======================================================
//  Structural coding
//=======================================================
// From Qsys

Computer_System The_System (
	////////////////////////////////////
	// FPGA Side
	////////////////////////////////////
	.vga_pio_locked_export			(vga_pll_lock),           //       vga_pio_locked.export
	.vga_pio_outclk0_clk				(vga_pll),              //      vga_pio_outclk0.clk
	.m10k_pll_locked_export			(M10k_pll_locked),          //      m10k_pll_locked.export
	.m10k_pll_outclk0_clk			(M10k_pll),            //     m10k_pll_outclk0.clk

	// Global signals
	.system_pll_ref_clk_clk					(CLOCK_50),
	.system_pll_ref_reset_reset			(1'b0),
	
	////////////////////////////////////
	// HPS Side
	////////////////////////////////////
	// DDR3 SDRAM
	.memory_mem_a			(HPS_DDR3_ADDR),
	.memory_mem_ba			(HPS_DDR3_BA),
	.memory_mem_ck			(HPS_DDR3_CK_P),
	.memory_mem_ck_n		(HPS_DDR3_CK_N),
	.memory_mem_cke		(HPS_DDR3_CKE),
	.memory_mem_cs_n		(HPS_DDR3_CS_N),
	.memory_mem_ras_n		(HPS_DDR3_RAS_N),
	.memory_mem_cas_n		(HPS_DDR3_CAS_N),
	.memory_mem_we_n		(HPS_DDR3_WE_N),
	.memory_mem_reset_n	(HPS_DDR3_RESET_N),
	.memory_mem_dq			(HPS_DDR3_DQ),
	.memory_mem_dqs		(HPS_DDR3_DQS_P),
	.memory_mem_dqs_n		(HPS_DDR3_DQS_N),
	.memory_mem_odt		(HPS_DDR3_ODT),
	.memory_mem_dm			(HPS_DDR3_DM),
	.memory_oct_rzqin		(HPS_DDR3_RZQ),
		  
	// Ethernet
	.hps_io_hps_io_gpio_inst_GPIO35	(HPS_ENET_INT_N),
	.hps_io_hps_io_emac1_inst_TX_CLK	(HPS_ENET_GTX_CLK),
	.hps_io_hps_io_emac1_inst_TXD0	(HPS_ENET_TX_DATA[0]),
	.hps_io_hps_io_emac1_inst_TXD1	(HPS_ENET_TX_DATA[1]),
	.hps_io_hps_io_emac1_inst_TXD2	(HPS_ENET_TX_DATA[2]),
	.hps_io_hps_io_emac1_inst_TXD3	(HPS_ENET_TX_DATA[3]),
	.hps_io_hps_io_emac1_inst_RXD0	(HPS_ENET_RX_DATA[0]),
	.hps_io_hps_io_emac1_inst_MDIO	(HPS_ENET_MDIO),
	.hps_io_hps_io_emac1_inst_MDC		(HPS_ENET_MDC),
	.hps_io_hps_io_emac1_inst_RX_CTL	(HPS_ENET_RX_DV),
	.hps_io_hps_io_emac1_inst_TX_CTL	(HPS_ENET_TX_EN),
	.hps_io_hps_io_emac1_inst_RX_CLK	(HPS_ENET_RX_CLK),
	.hps_io_hps_io_emac1_inst_RXD1	(HPS_ENET_RX_DATA[1]),
	.hps_io_hps_io_emac1_inst_RXD2	(HPS_ENET_RX_DATA[2]),
	.hps_io_hps_io_emac1_inst_RXD3	(HPS_ENET_RX_DATA[3]),

	// Flash
	.hps_io_hps_io_qspi_inst_IO0	(HPS_FLASH_DATA[0]),
	.hps_io_hps_io_qspi_inst_IO1	(HPS_FLASH_DATA[1]),
	.hps_io_hps_io_qspi_inst_IO2	(HPS_FLASH_DATA[2]),
	.hps_io_hps_io_qspi_inst_IO3	(HPS_FLASH_DATA[3]),
	.hps_io_hps_io_qspi_inst_SS0	(HPS_FLASH_NCSO),
	.hps_io_hps_io_qspi_inst_CLK	(HPS_FLASH_DCLK),

	// Accelerometer
	.hps_io_hps_io_gpio_inst_GPIO61	(HPS_GSENSOR_INT),

	//.adc_sclk                        (ADC_SCLK),
	//.adc_cs_n                        (ADC_CS_N),
	//.adc_dout                        (ADC_DOUT),
	//.adc_din                         (ADC_DIN),

	// General Purpose I/O
	.hps_io_hps_io_gpio_inst_GPIO40	(HPS_GPIO[0]),
	.hps_io_hps_io_gpio_inst_GPIO41	(HPS_GPIO[1]),

	// I2C
	.hps_io_hps_io_gpio_inst_GPIO48	(HPS_I2C_CONTROL),
	.hps_io_hps_io_i2c0_inst_SDA		(HPS_I2C1_SDAT),
	.hps_io_hps_io_i2c0_inst_SCL		(HPS_I2C1_SCLK),
	.hps_io_hps_io_i2c1_inst_SDA		(HPS_I2C2_SDAT),
	.hps_io_hps_io_i2c1_inst_SCL		(HPS_I2C2_SCLK),

	// Pushbutton
	.hps_io_hps_io_gpio_inst_GPIO54	(HPS_KEY),

	// LED
	.hps_io_hps_io_gpio_inst_GPIO53	(HPS_LED),

	// SD Card
	.hps_io_hps_io_sdio_inst_CMD	(HPS_SD_CMD),
	.hps_io_hps_io_sdio_inst_D0	(HPS_SD_DATA[0]),
	.hps_io_hps_io_sdio_inst_D1	(HPS_SD_DATA[1]),
	.hps_io_hps_io_sdio_inst_CLK	(HPS_SD_CLK),
	.hps_io_hps_io_sdio_inst_D2	(HPS_SD_DATA[2]),
	.hps_io_hps_io_sdio_inst_D3	(HPS_SD_DATA[3]),

	// SPI
	.hps_io_hps_io_spim1_inst_CLK		(HPS_SPIM_CLK),
	.hps_io_hps_io_spim1_inst_MOSI	(HPS_SPIM_MOSI),
	.hps_io_hps_io_spim1_inst_MISO	(HPS_SPIM_MISO),
	.hps_io_hps_io_spim1_inst_SS0		(HPS_SPIM_SS),

	// UART
	.hps_io_hps_io_uart0_inst_RX	(HPS_UART_RX),
	.hps_io_hps_io_uart0_inst_TX	(HPS_UART_TX),

	// USB
	.hps_io_hps_io_gpio_inst_GPIO09	(HPS_CONV_USB_N),
	.hps_io_hps_io_usb1_inst_D0		(HPS_USB_DATA[0]),
	.hps_io_hps_io_usb1_inst_D1		(HPS_USB_DATA[1]),
	.hps_io_hps_io_usb1_inst_D2		(HPS_USB_DATA[2]),
	.hps_io_hps_io_usb1_inst_D3		(HPS_USB_DATA[3]),
	.hps_io_hps_io_usb1_inst_D4		(HPS_USB_DATA[4]),
	.hps_io_hps_io_usb1_inst_D5		(HPS_USB_DATA[5]),
	.hps_io_hps_io_usb1_inst_D6		(HPS_USB_DATA[6]),
	.hps_io_hps_io_usb1_inst_D7		(HPS_USB_DATA[7]),
	.hps_io_hps_io_usb1_inst_CLK		(HPS_USB_CLKOUT),
	.hps_io_hps_io_usb1_inst_STP		(HPS_USB_STP),
	.hps_io_hps_io_usb1_inst_DIR		(HPS_USB_DIR),
	.hps_io_hps_io_usb1_inst_NXT		(HPS_USB_NXT),
	
	// counting render time
	.counter_external_connection_export(counter_external_connection_export),
	
	// wires for ci/cr increment/zoom and pio reset
	.pio_ci_init_external_connection_export(pio_ci_init_external_connection_export),
	.pio_cr_init_external_connection_export(pio_cr_init_external_connection_export),
	.pio_zoom_ci_external_connection_export(pio_zoom_ci_external_connection_export),
	.pio_zoom_cr_external_connection_export(pio_zoom_cr_external_connection_export),
	.pio_reset_external_connection_export(pio_reset_external_connection_export),
	
	// wire for max iterations
	.pio_max_iter_external_connection_export(pio_max_iter_external_connection_export)
);
endmodule // end top level

// color write data module
module color_write(clk, counter, max_iterations, write_data_out);
	input clk;
	input [11:0] counter, max_iterations;
	output [7:0] write_data_out;

	reg [7:0] write_data;

	always@(posedge clk) begin
		if (counter >= max_iterations) begin
		  write_data <= 8'b_000_000_00 ; // black
		end
		else if (counter >= (max_iterations >>> 1)) begin
		  write_data <= 8'b_011_001_00 ; 
		end
		else if (counter >= (max_iterations >>> 2)) begin
		  write_data <= 8'b_011_001_00 ;
		end
		else if (counter >= (max_iterations >>> 3)) begin
		  write_data <= 8'b_101_010_01 ;
		end
		else if (counter >= (max_iterations >>> 4)) begin
		  write_data <= 8'b_011_001_01 ;
		end
		else if (counter >= (max_iterations >>> 5)) begin
		  write_data <= 8'b_001_001_01 ;
		end
		else if (counter >= (max_iterations >>> 6)) begin
		  write_data <= 8'b_011_010_10 ;
		end
		else if (counter >= (max_iterations >>> 7)) begin
		  write_data <= 8'b_010_100_10 ;
		end
		else if (counter >= (max_iterations >>> 8)) begin
		  write_data <= 8'b_010_100_10 ; 
		end
		else begin
		  write_data <= 8'b_010_100_10 ;
		end
	end
	
	assign write_data_out = write_data;
endmodule

/*
// Key debouncing logic
module key_debouncing(clk,button_in,button_state);
	input clk, button_in;
	output [1:0] button_state;

	reg possible_button_press;
	reg [1:0] track_button;
	
	always @(posedge clk) begin
		if (track_button == 2'd0) begin //not pressed
			if (~button_in) begin
				track_button <= 2'd1;
				possible_button_press <= (~button_in);
			end
		end
		else if (track_button == 2'd1) begin //maybe pressed
			if ((~button_in) && possible_button_press) begin
				track_button <= 2'd2;
			end
			else begin
				track_button <= 2'd0;
			end
		end
		else if (track_button == 2'd2) begin //pressed
			if (button_in && possible_button_press) begin
				track_button <= 2'd3;
			end
			else begin
				track_button <= 2'd2;
			end
		end
		else if (track_button == 2'd3) begin //maybe not pressed
			if ((~button_in) && possible_button_press) begin
				track_button <= 2'd2;
			end
			else begin
				track_button <= 2'd0;
			end
		end
	end
	
	assign button_state = track_button;
endmodule
*/

// Declaration of module, include width and signedness of each input/output
module vga_driver (
	input wire clock,
	input wire reset,
	input [7:0] color_in,
	output [9:0] next_x,
	output [9:0] next_y,
	output wire hsync,
	output wire vsync,
	output [7:0] red,
	output [7:0] green,
	output [7:0] blue,
	output sync,
	output clk,
	output blank
);
	
	// Horizontal parameters (measured in clock cycles)
	parameter [9:0] H_ACTIVE  	=  10'd_639 ;
	parameter [9:0] H_FRONT 	=  10'd_15 ;
	parameter [9:0] H_PULSE		=  10'd_95 ;
	parameter [9:0] H_BACK 		=  10'd_47 ;

	// Vertical parameters (measured in lines)
	parameter [9:0] V_ACTIVE  	=  10'd_479 ;
	parameter [9:0] V_FRONT 	=  10'd_9 ;
	parameter [9:0] V_PULSE		=  10'd_1 ;
	parameter [9:0] V_BACK 		=  10'd_32 ;

//	// Horizontal parameters (measured in clock cycles)
//	parameter [9:0] H_ACTIVE  	=  10'd_9 ;
//	parameter [9:0] H_FRONT 	=  10'd_4 ;
//	parameter [9:0] H_PULSE		=  10'd_4 ;
//	parameter [9:0] H_BACK 		=  10'd_4 ;
//	parameter [9:0] H_TOTAL 	=  10'd_799 ;
//
//	// Vertical parameters (measured in lines)
//	parameter [9:0] V_ACTIVE  	=  10'd_1 ;
//	parameter [9:0] V_FRONT 	=  10'd_1 ;
//	parameter [9:0] V_PULSE		=  10'd_1 ;
//	parameter [9:0] V_BACK 		=  10'd_1 ;

	// Parameters for readability
	parameter 	LOW 	= 1'b_0 ;
	parameter 	HIGH	= 1'b_1 ;

	// States (more readable)
	parameter 	[7:0]	H_ACTIVE_STATE 		= 8'd_0 ;
	parameter 	[7:0] 	H_FRONT_STATE		= 8'd_1 ;
	parameter 	[7:0] 	H_PULSE_STATE 		= 8'd_2 ;
	parameter 	[7:0] 	H_BACK_STATE 		= 8'd_3 ;

	parameter 	[7:0]	V_ACTIVE_STATE 		= 8'd_0 ;
	parameter 	[7:0] 	V_FRONT_STATE		= 8'd_1 ;
	parameter 	[7:0] 	V_PULSE_STATE 		= 8'd_2 ;
	parameter 	[7:0] 	V_BACK_STATE 		= 8'd_3 ;

	// Clocked registers
	reg 		hysnc_reg ;
	reg 		vsync_reg ;
	reg 	[7:0]	red_reg ;
	reg 	[7:0]	green_reg ;
	reg 	[7:0]	blue_reg ;
	reg 		line_done ;

	// Control registers
	reg 	[9:0] 	h_counter ;
	reg 	[9:0] 	v_counter ;

	reg 	[7:0]	h_state ;
	reg 	[7:0]	v_state ;

	// State machine
	always@(posedge clock) begin
		// At reset . . .
  		if (reset) begin
			// Zero the counters
			h_counter 	<= 10'd_0 ;
			v_counter 	<= 10'd_0 ;
			// States to ACTIVE
			h_state 	<= H_ACTIVE_STATE  ;
			v_state 	<= V_ACTIVE_STATE  ;
			// Deassert line done
			line_done 	<= LOW ;
  		end
  		else begin
			//////////////////////////////////////////////////////////////////////////
			///////////////////////// HORIZONTAL /////////////////////////////////////
			//////////////////////////////////////////////////////////////////////////
			if (h_state == H_ACTIVE_STATE) begin
				// Iterate horizontal counter, zero at end of ACTIVE mode
				h_counter <= (h_counter==H_ACTIVE)?10'd_0:(h_counter + 10'd_1) ;
				// Set hsync
				hysnc_reg <= HIGH ;
				// Deassert line done
				line_done <= LOW ;
				// State transition
				h_state <= (h_counter == H_ACTIVE)?H_FRONT_STATE:H_ACTIVE_STATE ;
			end
			// Assert done flag, wait here for reset
			if (h_state == H_FRONT_STATE) begin
				// Iterate horizontal counter, zero at end of H_FRONT mode
				h_counter <= (h_counter==H_FRONT)?10'd_0:(h_counter + 10'd_1) ;
				// Set hsync
				hysnc_reg <= HIGH ;
				// State transition
				h_state <= (h_counter == H_FRONT)?H_PULSE_STATE:H_FRONT_STATE ;
			end
			if (h_state == H_PULSE_STATE) begin
				// Iterate horizontal counter, zero at end of H_FRONT mode
				h_counter <= (h_counter==H_PULSE)?10'd_0:(h_counter + 10'd_1) ;
				// Set hsync
				hysnc_reg <= LOW ;
				// State transition
				h_state <= (h_counter == H_PULSE)?H_BACK_STATE:H_PULSE_STATE ;
			end
			if (h_state == H_BACK_STATE) begin
				// Iterate horizontal counter, zero at end of H_FRONT mode
				h_counter <= (h_counter==H_BACK)?10'd_0:(h_counter + 10'd_1) ;
				// Set hsync
				hysnc_reg <= HIGH ;
				// State transition
				h_state <= (h_counter == H_BACK)?H_ACTIVE_STATE:H_BACK_STATE ;
				// Signal line complete at state transition (offset by 1 for synchronous state transition)
				line_done <= (h_counter == (H_BACK-1))?HIGH:LOW ;
			end
			//////////////////////////////////////////////////////////////////////////
			///////////////////////// VERTICAL ///////////////////////////////////////
			//////////////////////////////////////////////////////////////////////////
			if (v_state == V_ACTIVE_STATE) begin
				// increment vertical counter at end of line, zero on state transition
				v_counter <= (line_done==HIGH)?((v_counter==V_ACTIVE)?10'd_0:(v_counter + 10'd_1)):v_counter ;
				// set vsync in active mode
				vsync_reg <= HIGH ;
				// state transition - only on end of lines
				v_state <= (line_done==HIGH)?((v_counter==V_ACTIVE)?V_FRONT_STATE:V_ACTIVE_STATE):V_ACTIVE_STATE ;
			end
			if (v_state == V_FRONT_STATE) begin
				// increment vertical counter at end of line, zero on state transition
				v_counter <= (line_done==HIGH)?((v_counter==V_FRONT)?10'd_0:(v_counter + 10'd_1)):v_counter ;
				// set vsync in front porch
				vsync_reg <= HIGH ;
				// state transition
				v_state <= (line_done==HIGH)?((v_counter==V_FRONT)?V_PULSE_STATE:V_FRONT_STATE):V_FRONT_STATE ;
			end
			if (v_state == V_PULSE_STATE) begin
				// increment vertical counter at end of line, zero on state transition
				v_counter <= (line_done==HIGH)?((v_counter==V_PULSE)?10'd_0:(v_counter + 10'd_1)):v_counter ;
				// clear vsync in pulse
				vsync_reg <= LOW ;
				// state transition
				v_state <= (line_done==HIGH)?((v_counter==V_PULSE)?V_BACK_STATE:V_PULSE_STATE):V_PULSE_STATE ;
			end
			if (v_state == V_BACK_STATE) begin
				// increment vertical counter at end of line, zero on state transition
				v_counter <= (line_done==HIGH)?((v_counter==V_BACK)?10'd_0:(v_counter + 10'd_1)):v_counter ;
				// set vsync in back porch
				vsync_reg <= HIGH ;
				// state transition
				v_state <= (line_done==HIGH)?((v_counter==V_BACK)?V_ACTIVE_STATE:V_BACK_STATE):V_BACK_STATE ;
			end

			//////////////////////////////////////////////////////////////////////////
			//////////////////////////////// COLOR OUT ///////////////////////////////
			//////////////////////////////////////////////////////////////////////////
			red_reg 		<= (h_state==H_ACTIVE_STATE)?((v_state==V_ACTIVE_STATE)?{color_in[7:5],5'd_0}:8'd_0):8'd_0 ;
			green_reg 	<= (h_state==H_ACTIVE_STATE)?((v_state==V_ACTIVE_STATE)?{color_in[4:2],5'd_0}:8'd_0):8'd_0 ;
			blue_reg 	<= (h_state==H_ACTIVE_STATE)?((v_state==V_ACTIVE_STATE)?{color_in[1:0],6'd_0}:8'd_0):8'd_0 ;
			
 	 	end
	end
	// Assign output values
	assign hsync = hysnc_reg ;
	assign vsync = vsync_reg ;
	assign red = red_reg ;
	assign green = green_reg ;
	assign blue = blue_reg ;
	assign clk = clock ;
	assign sync = 1'b_0 ;
	assign blank = hysnc_reg & vsync_reg ;
	// The x/y coordinates that should be available on the NEXT cycle
	assign next_x = (h_state==H_ACTIVE_STATE)?h_counter:10'd_0 ;
	assign next_y = (v_state==V_ACTIVE_STATE)?v_counter:10'd_0 ;

endmodule

//////////////////////////////////////////////////////////////
////////////	Mandelbrot Set Visualizer	    //////////////
//////////////////////////////////////////////////////////////

module mandelbrot (clock, reset, x_coord_init, y_coord_init, step_size_cr, step_size_ci, c_i_init, c_r_init, max_iter, out, write_en, write_addr, done, time_flag, time_counter);
   input clock, reset;
	input [9:0] x_coord_init, y_coord_init;
	input signed [26:0] c_i_init, c_r_init;
	input signed [26:0] step_size_cr, step_size_ci;
	input [11:0] max_iter;
	output [11:0] out;
	output [18:0] write_addr;
	output write_en;
	output done;
	output time_flag;
	output [31:0] time_counter;
	
	reg t_flag;
	reg [31:0] running_counter, t_counter;
	
	reg write_enable;
	reg [1:0] state;
	reg [9:0] x_coord, y_coord;
	reg signed [26:0] ci, cr;
	reg [18:0] write_address;
   reg signed [26:0] z_r, z_i;
   reg [11:0] temp_iter;
   wire signed [26:0] zr_sq, zi_sq, zr_zi;
   wire signed [26:0] zr_temp, zi_temp;
	wire [26:0] zr_abs, zi_abs;

    // clocked
    always @(posedge clock) begin
		 if (reset == 1) begin
			z_r <= 0;
			z_i <= 0;
			x_coord <= x_coord_init;
			y_coord <= y_coord_init;
			temp_iter <= 0;
			ci <= c_i_init;
			cr <= c_r_init;
			state <= 2'd0;
			t_flag <= 1'd0;
			running_counter <= 32'd0; 
			t_counter <= 32'd0;
			write_enable <= 1'd0;
			write_address <= 19'd0;
		
		 end
		 else begin
			if (state == 0) begin
					z_r <= 0;
					z_i <= 0;
					temp_iter <= 0;
					state <= 1;
					write_enable <= 1'd0;
			end
			else if (state == 1) begin
				if (~done) begin
					z_r <= zr_temp;
					z_i <= zi_temp;
					temp_iter <= temp_iter + 1;
					state <= 1;
				end
				else begin
					state <= 2;
				end
			end
			else if (state == 2) begin
				write_enable <= 1'd1;
				write_address <= (19'd_40 * y_coord) + (x_coord >> 4);
				x_coord <= (x_coord==10'd_624 + x_coord_init) ? (x_coord_init) : (x_coord + 10'd_16) ;
				y_coord <= (x_coord==10'd_624 + x_coord_init) ? ((y_coord==10'd_479) ? 10'd_0 : (y_coord+10'd_1)) : y_coord ;
				cr <= (x_coord==10'd_624 + x_coord_init) ? (c_r_init) : (cr + step_size_cr); //{4'b0000,23'b00000010011001100110010} // x
				ci <= (x_coord==10'd_624 + x_coord_init) ? ((y_coord==10'd_479) ? (c_i_init): (ci - step_size_ci)) : ci ; // y
				state <= 0;
				t_flag <= ((x_coord==10'd_624 + x_coord_init) && (y_coord==10'd_479)) ? 1 : 0;
			end
//			running_counter <= (t_flag == 0) ? (running_counter + 32'd1) : running_counter;
			if (t_flag != 1) begin
//				t_counter <= running_counter;
				running_counter <= (running_counter + 32'd1);
//	         t_flag <= 0;
//				running_counter <= 0;
			end
			else begin
				running_counter <= 0;
			end
		end
    end
   
    // signed mults
    signed_mult zrSq (.out(zr_sq), .a(z_r), .b(z_r));
    signed_mult ziSq (.out(zi_sq), .a(z_i), .b(z_i));
    signed_mult twoZrZi (.out(zr_zi), .a(z_r), .b(z_i));

    // combinational
	 assign time_flag = t_flag;
	 assign time_counter = running_counter;
    assign zr_temp = zr_sq - zi_sq + cr;
    assign zi_temp = (zr_zi <<< 1) + ci;
	 assign zr_abs = (z_r[26] == 1) ? (~z_r + 1) : (z_r);  
	 assign zi_abs = (z_i[26] == 1) ? (~z_i + 1) : (z_i);  
    assign done = (zr_abs > {4'd2, 23'd0}) || (zi_abs > {4'd2, 23'd0}) || ((zr_sq + zi_sq) > {4'd4, 23'd0}) || (temp_iter >= max_iter); 
	 assign out = temp_iter;
	 assign write_en = write_enable;
	 assign write_addr = write_address;
endmodule

//////////////////////////////////////////////////
//// signed mult of 4.23 format 2'comp////////////
//////////////////////////////////////////////////
module signed_mult (out, a, b);
	output 	signed  [26:0]	out;
	input 	signed	[26:0] 	a;
	input 	signed	[26:0] 	b;
    
	// intermediate full bit length
	wire 	signed	[53:0]	mult_out;
	assign mult_out = a * b;
    
	// select bits for 4.23 fixed point
	assign out = {mult_out[53], mult_out[48:23]};
endmodule


//============================================================
// M10K module for testing
//============================================================
// See example 12-16 in 
// http://people.ece.cornell.edu/land/courses/ece5760/DE1_SOC/HDL_style_qts_qii51007.pdf
//============================================================

module M10K_1000_8( 
    output reg [7:0] q,
    input [7:0] d,
    input [18:0] write_address, read_address,
    input we, clk
);
	 // force M10K ram style
	 // 307200 words of 8 bits
	 //307200
    reg [7:0] mem [19200:0]  /* synthesis ramstyle = "no_rw_check, M10K" */;
	 
    always @ (posedge clk) begin
        if (we) begin
            mem[write_address] <= d;
		  end
		  
        q <= mem[read_address]; // q doesn't get d in this clock cycle
    end
endmodule
